package shared_pkg;
    typedef enum  {OR,XOR,ADD,MULT,SHIFT,ROTATE,INVALID_6,INVALID_7} opcode_e;
    localparam MAXPOS = 3 , MAXNEG = -4 , ZERO = 0;
endpackage